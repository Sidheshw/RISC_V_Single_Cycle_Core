module PC_adder(a , b ,c);

input [31:0] a , b ;
input [31:0] c;

assign c=a+b;


endmodule